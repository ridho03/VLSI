magic
tech sky130A
magscale 1 2
timestamp 1729218614
<< psubdiff >>
rect 2801 1486 2861 1520
rect 3920 1486 3980 1520
rect 2801 1460 2835 1486
rect 3946 1460 3980 1486
rect 2801 -7 2835 19
rect 3946 -7 3980 19
rect 2801 -41 2861 -7
rect 3920 -41 3980 -7
<< psubdiffcont >>
rect 2861 1486 3920 1520
rect 2801 19 2835 1460
rect 3946 19 3980 1460
rect 2861 -41 3920 -7
<< poly >>
rect 2920 1334 3012 1350
rect 2920 1300 2936 1334
rect 2970 1300 3012 1334
rect 2920 1284 3012 1300
rect 2982 1250 3012 1284
rect 3738 1330 3830 1346
rect 3738 1296 3780 1330
rect 3814 1296 3830 1330
rect 3738 1280 3830 1296
rect 3738 1246 3768 1280
rect 3070 666 3680 778
rect 2982 150 3012 184
rect 2920 134 3012 150
rect 2920 100 2936 134
rect 2970 100 3012 134
rect 2920 84 3012 100
rect 3738 145 3768 179
rect 3738 129 3830 145
rect 3738 95 3780 129
rect 3814 95 3830 129
rect 3738 79 3830 95
<< polycont >>
rect 2936 1300 2970 1334
rect 3780 1296 3814 1330
rect 2936 100 2970 134
rect 3780 95 3814 129
<< locali >>
rect 2801 1486 2861 1520
rect 3920 1486 3980 1520
rect 2801 1460 2835 1486
rect 3946 1460 3980 1486
rect 2920 1300 2936 1334
rect 2970 1300 2986 1334
rect 2936 1250 2970 1300
rect 3764 1296 3780 1330
rect 3814 1296 3830 1330
rect 3780 1246 3814 1296
rect 2936 134 2970 184
rect 2920 100 2936 134
rect 2970 100 2986 134
rect 3780 129 3814 179
rect 3764 95 3780 129
rect 3814 95 3830 129
rect 2801 -7 2835 19
rect 3946 -7 3980 19
rect 2801 -41 2861 -7
rect 3920 -41 3980 -7
<< viali >>
rect 3282 1486 3316 1520
rect 2936 1300 2970 1334
rect 3780 1296 3814 1330
rect 2936 100 2970 134
rect 3780 95 3814 129
rect 3433 -41 3470 -7
<< metal1 >>
rect 3269 1477 3279 1529
rect 3331 1477 3341 1529
rect 2924 1334 2982 1340
rect 2924 1300 2936 1334
rect 2970 1300 2982 1334
rect 2924 1294 2982 1300
rect 3768 1330 3826 1336
rect 3768 1296 3780 1330
rect 3814 1296 3826 1330
rect 2930 1250 2976 1294
rect 3768 1290 3826 1296
rect 3774 1251 3820 1290
rect 2924 850 3070 1249
rect 3680 1238 3826 1251
rect 3263 862 3273 1238
rect 3325 862 3335 1238
rect 3415 862 3425 1238
rect 3477 862 3487 1238
rect 3673 862 3683 1238
rect 3735 862 3826 1238
rect 3680 852 3826 862
rect 3024 812 3058 850
rect 3024 778 3108 812
rect 3238 778 3391 812
rect 3357 650 3391 778
rect 3357 616 3517 650
rect 3648 610 3726 656
rect 2924 566 3077 579
rect 3692 578 3726 610
rect 2924 190 3015 566
rect 3067 190 3077 566
rect 3263 190 3273 566
rect 3325 190 3335 566
rect 3415 190 3425 566
rect 3477 190 3487 566
rect 2924 179 3077 190
rect 3680 179 3826 578
rect 2930 140 2976 179
rect 2924 134 2982 140
rect 3774 135 3820 179
rect 2924 100 2936 134
rect 2970 100 2982 134
rect 2924 94 2982 100
rect 3768 129 3826 135
rect 3768 95 3780 129
rect 3814 95 3826 129
rect 3768 89 3826 95
rect 3416 -50 3426 2
rect 3478 -50 3488 2
<< via1 >>
rect 3279 1520 3331 1529
rect 3279 1486 3282 1520
rect 3282 1486 3316 1520
rect 3316 1486 3331 1520
rect 3279 1477 3331 1486
rect 3273 862 3325 1238
rect 3425 862 3477 1238
rect 3683 862 3735 1238
rect 3015 190 3067 566
rect 3273 190 3325 566
rect 3425 190 3477 566
rect 3426 -7 3478 2
rect 3426 -41 3433 -7
rect 3433 -41 3470 -7
rect 3470 -41 3478 -7
rect 3426 -50 3478 -41
<< metal2 >>
rect 3277 1531 3333 1541
rect 3277 1465 3333 1475
rect 3271 1238 3327 1248
rect 3271 852 3327 862
rect 3423 1238 3479 1248
rect 3683 1238 3735 1248
rect 3423 852 3479 862
rect 3673 862 3683 884
rect 3735 862 3745 884
rect 3673 818 3745 862
rect 3339 746 3745 818
rect 3339 681 3411 746
rect 3005 609 3411 681
rect 3005 566 3077 609
rect 3005 553 3015 566
rect 3067 553 3077 566
rect 3271 566 3327 576
rect 3015 180 3067 190
rect 3271 180 3327 190
rect 3423 566 3479 576
rect 3423 180 3479 190
rect 3424 4 3480 14
rect 3424 -62 3480 -52
<< via2 >>
rect 3277 1529 3333 1531
rect 3277 1477 3279 1529
rect 3279 1477 3331 1529
rect 3331 1477 3333 1529
rect 3277 1475 3333 1477
rect 3271 862 3273 1238
rect 3273 862 3325 1238
rect 3325 862 3327 1238
rect 3423 862 3425 1238
rect 3425 862 3477 1238
rect 3477 862 3479 1238
rect 3271 190 3273 566
rect 3273 190 3325 566
rect 3325 190 3327 566
rect 3423 190 3425 566
rect 3425 190 3477 566
rect 3477 190 3479 566
rect 3424 2 3480 4
rect 3424 -50 3426 2
rect 3426 -50 3478 2
rect 3478 -50 3480 2
rect 3424 -52 3480 -50
<< metal3 >>
rect 3252 1536 3357 1550
rect 3252 1472 3273 1536
rect 3337 1472 3357 1536
rect 3252 1456 3357 1472
rect 3261 1238 3337 1243
rect 3413 1238 3489 1243
rect 3257 862 3267 1238
rect 3331 862 3341 1238
rect 3413 862 3423 1238
rect 3479 862 3489 1238
rect 3261 857 3337 862
rect 3413 742 3489 862
rect 3261 666 3489 742
rect 3261 566 3337 666
rect 3413 566 3489 571
rect 3261 190 3271 566
rect 3327 190 3337 566
rect 3409 190 3419 566
rect 3483 190 3493 566
rect 3261 185 3337 190
rect 3413 185 3489 190
rect 3396 8 3505 24
rect 3396 -56 3420 8
rect 3484 -56 3505 8
rect 3396 -71 3505 -56
<< via3 >>
rect 3273 1531 3337 1536
rect 3273 1475 3277 1531
rect 3277 1475 3333 1531
rect 3333 1475 3337 1531
rect 3273 1472 3337 1475
rect 3267 862 3271 1238
rect 3271 862 3327 1238
rect 3327 862 3331 1238
rect 3419 190 3423 566
rect 3423 190 3479 566
rect 3479 190 3483 566
rect 3420 4 3484 8
rect 3420 -52 3424 4
rect 3424 -52 3480 4
rect 3480 -52 3484 4
rect 3420 -56 3484 -52
<< metal4 >>
rect 3272 1536 3338 1537
rect 3272 1494 3273 1536
rect 3257 1472 3273 1494
rect 3337 1494 3338 1536
rect 3337 1472 3341 1494
rect 3257 1238 3341 1472
rect 3257 1229 3267 1238
rect 3266 878 3267 1229
rect 3257 862 3267 878
rect 3331 1229 3341 1238
rect 3331 878 3332 1229
rect 3331 862 3341 878
rect 3257 756 3341 862
rect 3257 672 3492 756
rect 3408 566 3492 672
rect 3408 556 3419 566
rect 3418 201 3419 556
rect 3407 190 3419 201
rect 3483 556 3492 566
rect 3483 201 3484 556
rect 3483 190 3492 201
rect 3407 8 3492 190
rect 3407 -15 3420 8
rect 3419 -56 3420 -15
rect 3484 -15 3492 8
rect 3484 -56 3485 -15
rect 3419 -57 3485 -56
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_0
timestamp 1729218115
transform 1 0 3170 0 1 1050
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_1
timestamp 1729218115
transform 1 0 3580 0 1 1050
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_2
timestamp 1729218115
transform 1 0 3170 0 1 378
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_3
timestamp 1729218115
transform 1 0 3580 0 1 378
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_4
timestamp 1729168343
transform 1 0 2997 0 1 378
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_5
timestamp 1729168343
transform 1 0 3753 0 1 378
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_6
timestamp 1729168343
transform 1 0 2997 0 1 1050
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_7
timestamp 1729168343
transform 1 0 3753 0 1 1050
box -73 -226 73 226
<< labels >>
flabel metal4 3301 1370 3301 1370 0 FreeSans 640 0 0 0 gnd
port 0 nsew
flabel metal1 3034 804 3034 804 0 FreeSans 640 0 0 0 d3
port 1 nsew
flabel metal3 3456 824 3456 824 0 FreeSans 640 0 0 0 rs
port 2 nsew
flabel metal2 3717 804 3717 804 0 FreeSans 640 0 0 0 d4
port 3 nsew
<< end >>
