magic
tech sky130A
timestamp 1729184360
<< pwell >>
rect -148 -174 148 174
<< nmos >>
rect -50 -100 50 100
<< ndiff >>
rect -79 94 -50 100
rect -79 -94 -73 94
rect -56 -94 -50 94
rect -79 -100 -50 -94
rect 50 94 79 100
rect 50 -94 56 94
rect 73 -94 79 94
rect 50 -100 79 -94
<< ndiffc >>
rect -73 -94 -56 94
rect 56 -94 73 94
<< psubdiff >>
rect -130 139 -82 156
rect 82 139 130 156
rect -130 108 -113 139
rect 113 108 130 139
rect -130 -139 -113 -108
rect 113 -139 130 -108
rect -130 -156 -82 -139
rect 82 -156 130 -139
<< psubdiffcont >>
rect -82 139 82 156
rect -130 -108 -113 108
rect 113 -108 130 108
rect -82 -156 82 -139
<< poly >>
rect -50 100 50 113
rect -50 -113 50 -100
<< locali >>
rect -130 139 -82 156
rect 82 139 130 156
rect -130 108 -113 139
rect 113 108 130 139
rect -73 94 -56 102
rect -73 -102 -56 -94
rect 56 94 73 102
rect 56 -102 73 -94
rect -130 -139 -113 -108
rect 113 -139 130 -108
rect -130 -156 -82 -139
rect 82 -156 130 -139
<< viali >>
rect -73 -94 -56 94
rect 56 -94 73 94
<< metal1 >>
rect -76 94 -53 100
rect -76 -94 -73 94
rect -56 -94 -53 94
rect -76 -100 -53 -94
rect 53 94 76 100
rect 53 -94 56 94
rect 73 -94 76 94
rect 53 -100 76 -94
<< properties >>
string FIXED_BBOX -121 -147 121 147
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
