magic
tech sky130A
magscale 1 2
timestamp 1729158256
<< nwell >>
rect -232 53 767 2922
<< nsubdiff >>
rect -196 2852 -136 2886
rect 636 2852 731 2886
rect -196 2819 -162 2852
rect 697 2819 731 2852
rect -196 123 -162 149
rect 697 123 731 149
rect -196 89 -136 123
rect 636 89 731 123
<< nsubdiffcont >>
rect -136 2852 636 2886
rect -196 149 -162 2819
rect 697 149 731 2819
rect -136 89 636 123
<< poly >>
rect -111 2812 -19 2828
rect -111 2778 -95 2812
rect -61 2778 -19 2812
rect -111 2762 -19 2778
rect -49 2748 -19 2762
rect 555 2814 647 2830
rect 555 2780 597 2814
rect 631 2780 647 2814
rect 555 2764 647 2780
rect 555 2747 585 2764
rect -111 2114 -19 2130
rect 39 2129 239 2229
rect -111 2080 -95 2114
rect -61 2080 -19 2114
rect -111 2064 -19 2080
rect -49 2048 -19 2064
rect 555 2113 647 2129
rect 555 2079 597 2113
rect 631 2079 647 2113
rect 555 2063 647 2079
rect 555 2049 585 2063
rect 39 1435 497 1535
rect -49 899 -19 913
rect -111 883 -19 899
rect -111 849 -95 883
rect -61 849 -19 883
rect -111 833 -19 849
rect 555 903 585 917
rect 555 887 647 903
rect 555 853 597 887
rect 631 853 647 887
rect 296 739 497 841
rect 555 837 647 853
rect -50 211 -20 225
rect -112 195 -20 211
rect -112 161 -96 195
rect -62 161 -20 195
rect -112 145 -20 161
rect 554 211 584 225
rect 554 195 646 211
rect 554 161 596 195
rect 630 161 646 195
rect 554 145 646 161
<< polycont >>
rect -95 2778 -61 2812
rect 597 2780 631 2814
rect -95 2080 -61 2114
rect 597 2079 631 2113
rect -95 849 -61 883
rect 597 853 631 887
rect -96 161 -62 195
rect 596 161 630 195
<< locali >>
rect -196 2852 -136 2886
rect 636 2852 731 2886
rect -196 2819 -162 2852
rect 697 2819 731 2852
rect -111 2778 -95 2812
rect -61 2778 -45 2812
rect 581 2780 597 2814
rect 631 2780 647 2814
rect -95 2728 -61 2778
rect 597 2717 631 2780
rect -111 2080 -95 2114
rect -61 2080 -45 2114
rect -95 2025 -61 2080
rect 581 2079 597 2113
rect 631 2079 647 2113
rect 596 2014 631 2079
rect -95 883 -61 948
rect 597 887 631 958
rect -111 849 -95 883
rect -61 849 -45 883
rect 581 853 597 887
rect 631 853 647 887
rect -96 195 -62 262
rect 596 195 630 259
rect -112 161 -96 195
rect -62 161 -46 195
rect 580 161 596 195
rect 630 161 646 195
rect -196 123 -162 149
rect 697 123 731 149
rect -196 89 -136 123
rect 636 89 731 123
<< viali >>
rect 597 2852 631 2886
rect -95 2778 -61 2812
rect 597 2780 631 2814
rect -95 2080 -61 2114
rect 597 2079 631 2113
rect -95 849 -61 883
rect 597 853 631 887
rect -96 161 -62 195
rect 596 161 630 195
rect -96 89 -62 123
<< metal1 >>
rect 585 2886 643 2892
rect 585 2852 597 2886
rect 631 2852 643 2886
rect -107 2812 -49 2818
rect -107 2778 -95 2812
rect -61 2778 -49 2812
rect -107 2772 -49 2778
rect 585 2814 643 2852
rect 585 2780 597 2814
rect 631 2780 643 2814
rect 585 2774 643 2780
rect -101 2726 -55 2772
rect 592 2726 637 2774
rect -101 2714 33 2726
rect -114 2338 -104 2714
rect -52 2338 33 2714
rect -101 2326 33 2338
rect 244 2285 291 2726
rect 503 2345 637 2726
rect 502 2326 637 2345
rect 502 2285 549 2326
rect 244 2238 549 2285
rect -107 2114 -49 2120
rect -107 2080 -95 2114
rect -61 2080 -49 2114
rect -107 2074 -49 2080
rect -101 2032 -56 2074
rect -101 2020 27 2032
rect -101 1644 -16 2020
rect 36 1644 46 2020
rect -101 1632 27 1644
rect -7 1385 76 1419
rect -7 1338 27 1385
rect -101 1330 27 1338
rect -101 938 26 1330
rect -101 889 -55 938
rect -107 883 -49 889
rect -107 849 -95 883
rect -61 849 -49 883
rect -107 843 -49 849
rect 244 734 291 2238
rect 585 2113 643 2119
rect 585 2079 597 2113
rect 631 2079 643 2113
rect 585 2073 643 2079
rect 591 2032 637 2073
rect 503 1632 637 2032
rect 510 1584 543 1632
rect 462 1551 543 1584
rect 503 1326 630 1339
rect 490 950 500 1326
rect 552 958 630 1326
rect 552 950 637 958
rect 503 939 637 950
rect 591 893 637 939
rect 585 887 643 893
rect 585 853 597 887
rect 631 853 643 887
rect 585 847 643 853
rect -16 687 291 734
rect -16 642 31 687
rect -102 626 31 642
rect -102 242 32 626
rect 244 242 291 687
rect 508 630 632 642
rect 508 254 587 630
rect 639 254 649 630
rect -102 201 -57 242
rect 508 241 636 254
rect 591 201 636 241
rect -108 195 -50 201
rect -108 161 -96 195
rect -62 161 -50 195
rect -108 123 -50 161
rect 584 195 642 201
rect 584 161 596 195
rect 630 161 642 195
rect 584 155 642 161
rect -108 89 -96 123
rect -62 89 -50 123
rect -108 83 -50 89
<< via1 >>
rect -104 2338 -52 2714
rect -16 1644 36 2020
rect 500 950 552 1326
rect 587 254 639 630
<< metal2 >>
rect -104 2714 -52 2724
rect -104 2328 -52 2338
rect -95 2203 -61 2328
rect -95 2194 -38 2203
rect -95 2138 -94 2194
rect -95 2129 -38 2138
rect 575 2136 584 2196
rect 644 2136 653 2196
rect -95 831 -61 2129
rect -16 2020 36 2030
rect -16 1511 36 1644
rect -17 1459 551 1511
rect 500 1326 552 1459
rect 500 940 552 950
rect -108 822 -48 831
rect 596 829 631 2136
rect -108 753 -48 762
rect 572 820 631 829
rect 628 764 631 820
rect 572 755 631 764
rect 596 640 631 755
rect 587 630 639 640
rect 587 244 639 254
<< via2 >>
rect -94 2138 -38 2194
rect 584 2136 644 2196
rect -108 762 -48 822
rect 572 764 628 820
<< metal3 >>
rect -99 2196 -33 2199
rect 579 2196 649 2201
rect -99 2194 584 2196
rect -99 2138 -94 2194
rect -38 2138 584 2194
rect -99 2136 584 2138
rect 644 2136 649 2196
rect -99 2133 -33 2136
rect 579 2131 649 2136
rect -113 823 -43 827
rect 567 823 633 825
rect -113 822 633 823
rect -113 762 -108 822
rect -48 820 633 822
rect -48 764 572 820
rect 628 764 633 820
rect -48 762 633 764
rect -113 761 633 762
rect -113 757 -43 761
rect 567 759 633 761
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729135022
transform 1 0 -34 0 1 1832
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729135022
transform 1 0 -35 0 1 442
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729135022
transform 1 0 569 0 1 442
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729135022
transform 1 0 -34 0 1 1138
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729135022
transform 1 0 570 0 1 1138
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729135022
transform 1 0 570 0 1 1832
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729135022
transform 1 0 570 0 1 2526
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729135022
transform 1 0 -34 0 1 2526
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729135022
transform 1 0 268 0 1 2526
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729135022
transform 1 0 268 0 1 1832
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729135022
transform 1 0 268 0 1 1138
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729135022
transform 1 0 267 0 1 442
box -323 -300 323 300
<< labels >>
flabel metal2 617 1375 617 1375 0 FreeSans 1600 0 0 0 d5
port 3 nsew
flabel metal1 522 1586 522 1586 0 FreeSans 1600 0 0 0 d2
port 2 nsew
flabel metal2 14 1573 14 1573 0 FreeSans 1600 0 0 0 d1
port 1 nsew
flabel metal1 610 2840 610 2840 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
<< end >>
