magic
tech sky130A
magscale 1 2
timestamp 1729236880
<< nmos >>
rect -578 109 -418 309
rect -246 109 -86 309
rect 86 109 246 309
rect 418 109 578 309
rect -578 -309 -418 -109
rect -246 -309 -86 -109
rect 86 -309 246 -109
rect 418 -309 578 -109
<< ndiff >>
rect -636 297 -578 309
rect -636 121 -624 297
rect -590 121 -578 297
rect -636 109 -578 121
rect -418 297 -360 309
rect -418 121 -406 297
rect -372 121 -360 297
rect -418 109 -360 121
rect -304 297 -246 309
rect -304 121 -292 297
rect -258 121 -246 297
rect -304 109 -246 121
rect -86 297 -28 309
rect -86 121 -74 297
rect -40 121 -28 297
rect -86 109 -28 121
rect 28 297 86 309
rect 28 121 40 297
rect 74 121 86 297
rect 28 109 86 121
rect 246 297 304 309
rect 246 121 258 297
rect 292 121 304 297
rect 246 109 304 121
rect 360 297 418 309
rect 360 121 372 297
rect 406 121 418 297
rect 360 109 418 121
rect 578 297 636 309
rect 578 121 590 297
rect 624 121 636 297
rect 578 109 636 121
rect -636 -121 -578 -109
rect -636 -297 -624 -121
rect -590 -297 -578 -121
rect -636 -309 -578 -297
rect -418 -121 -360 -109
rect -418 -297 -406 -121
rect -372 -297 -360 -121
rect -418 -309 -360 -297
rect -304 -121 -246 -109
rect -304 -297 -292 -121
rect -258 -297 -246 -121
rect -304 -309 -246 -297
rect -86 -121 -28 -109
rect -86 -297 -74 -121
rect -40 -297 -28 -121
rect -86 -309 -28 -297
rect 28 -121 86 -109
rect 28 -297 40 -121
rect 74 -297 86 -121
rect 28 -309 86 -297
rect 246 -121 304 -109
rect 246 -297 258 -121
rect 292 -297 304 -121
rect 246 -309 304 -297
rect 360 -121 418 -109
rect 360 -297 372 -121
rect 406 -297 418 -121
rect 360 -309 418 -297
rect 578 -121 636 -109
rect 578 -297 590 -121
rect 624 -297 636 -121
rect 578 -309 636 -297
<< ndiffc >>
rect -624 121 -590 297
rect -406 121 -372 297
rect -292 121 -258 297
rect -74 121 -40 297
rect 40 121 74 297
rect 258 121 292 297
rect 372 121 406 297
rect 590 121 624 297
rect -624 -297 -590 -121
rect -406 -297 -372 -121
rect -292 -297 -258 -121
rect -74 -297 -40 -121
rect 40 -297 74 -121
rect 258 -297 292 -121
rect 372 -297 406 -121
rect 590 -297 624 -121
<< poly >>
rect -578 381 -418 397
rect -578 347 -562 381
rect -434 347 -418 381
rect -578 309 -418 347
rect -246 381 -86 397
rect -246 347 -230 381
rect -102 347 -86 381
rect -246 309 -86 347
rect 86 381 246 397
rect 86 347 102 381
rect 230 347 246 381
rect 86 309 246 347
rect 418 381 578 397
rect 418 347 434 381
rect 562 347 578 381
rect 418 309 578 347
rect -578 71 -418 109
rect -578 37 -562 71
rect -434 37 -418 71
rect -578 21 -418 37
rect -246 71 -86 109
rect -246 37 -230 71
rect -102 37 -86 71
rect -246 21 -86 37
rect 86 71 246 109
rect 86 37 102 71
rect 230 37 246 71
rect 86 21 246 37
rect 418 71 578 109
rect 418 37 434 71
rect 562 37 578 71
rect 418 21 578 37
rect -578 -37 -418 -21
rect -578 -71 -562 -37
rect -434 -71 -418 -37
rect -578 -109 -418 -71
rect -246 -37 -86 -21
rect -246 -71 -230 -37
rect -102 -71 -86 -37
rect -246 -109 -86 -71
rect 86 -37 246 -21
rect 86 -71 102 -37
rect 230 -71 246 -37
rect 86 -109 246 -71
rect 418 -37 578 -21
rect 418 -71 434 -37
rect 562 -71 578 -37
rect 418 -109 578 -71
rect -578 -347 -418 -309
rect -578 -381 -562 -347
rect -434 -381 -418 -347
rect -578 -397 -418 -381
rect -246 -347 -86 -309
rect -246 -381 -230 -347
rect -102 -381 -86 -347
rect -246 -397 -86 -381
rect 86 -347 246 -309
rect 86 -381 102 -347
rect 230 -381 246 -347
rect 86 -397 246 -381
rect 418 -347 578 -309
rect 418 -381 434 -347
rect 562 -381 578 -347
rect 418 -397 578 -381
<< polycont >>
rect -562 347 -434 381
rect -230 347 -102 381
rect 102 347 230 381
rect 434 347 562 381
rect -562 37 -434 71
rect -230 37 -102 71
rect 102 37 230 71
rect 434 37 562 71
rect -562 -71 -434 -37
rect -230 -71 -102 -37
rect 102 -71 230 -37
rect 434 -71 562 -37
rect -562 -381 -434 -347
rect -230 -381 -102 -347
rect 102 -381 230 -347
rect 434 -381 562 -347
<< locali >>
rect -578 347 -562 381
rect -434 347 -418 381
rect -246 347 -230 381
rect -102 347 -86 381
rect 86 347 102 381
rect 230 347 246 381
rect 418 347 434 381
rect 562 347 578 381
rect -624 297 -590 313
rect -624 105 -590 121
rect -406 297 -372 313
rect -406 105 -372 121
rect -292 297 -258 313
rect -292 105 -258 121
rect -74 297 -40 313
rect -74 105 -40 121
rect 40 297 74 313
rect 40 105 74 121
rect 258 297 292 313
rect 258 105 292 121
rect 372 297 406 313
rect 372 105 406 121
rect 590 297 624 313
rect 590 105 624 121
rect -578 37 -562 71
rect -434 37 -418 71
rect -246 37 -230 71
rect -102 37 -86 71
rect 86 37 102 71
rect 230 37 246 71
rect 418 37 434 71
rect 562 37 578 71
rect -578 -71 -562 -37
rect -434 -71 -418 -37
rect -246 -71 -230 -37
rect -102 -71 -86 -37
rect 86 -71 102 -37
rect 230 -71 246 -37
rect 418 -71 434 -37
rect 562 -71 578 -37
rect -624 -121 -590 -105
rect -624 -313 -590 -297
rect -406 -121 -372 -105
rect -406 -313 -372 -297
rect -292 -121 -258 -105
rect -292 -313 -258 -297
rect -74 -121 -40 -105
rect -74 -313 -40 -297
rect 40 -121 74 -105
rect 40 -313 74 -297
rect 258 -121 292 -105
rect 258 -313 292 -297
rect 372 -121 406 -105
rect 372 -313 406 -297
rect 590 -121 624 -105
rect 590 -313 624 -297
rect -578 -381 -562 -347
rect -434 -381 -418 -347
rect -246 -381 -230 -347
rect -102 -381 -86 -347
rect 86 -381 102 -347
rect 230 -381 246 -347
rect 418 -381 434 -347
rect 562 -381 578 -347
<< viali >>
rect -562 347 -434 381
rect -230 347 -102 381
rect 102 347 230 381
rect 434 347 562 381
rect -624 121 -590 297
rect -406 121 -372 297
rect -292 121 -258 297
rect -74 121 -40 297
rect 40 121 74 297
rect 258 121 292 297
rect 372 121 406 297
rect 590 121 624 297
rect -562 37 -434 71
rect -230 37 -102 71
rect 102 37 230 71
rect 434 37 562 71
rect -562 -71 -434 -37
rect -230 -71 -102 -37
rect 102 -71 230 -37
rect 434 -71 562 -37
rect -624 -297 -590 -121
rect -406 -297 -372 -121
rect -292 -297 -258 -121
rect -74 -297 -40 -121
rect 40 -297 74 -121
rect 258 -297 292 -121
rect 372 -297 406 -121
rect 590 -297 624 -121
rect -562 -381 -434 -347
rect -230 -381 -102 -347
rect 102 -381 230 -347
rect 434 -381 562 -347
<< metal1 >>
rect -574 381 -422 387
rect -574 347 -562 381
rect -434 347 -422 381
rect -574 341 -422 347
rect -242 381 -90 387
rect -242 347 -230 381
rect -102 347 -90 381
rect -242 341 -90 347
rect 90 381 242 387
rect 90 347 102 381
rect 230 347 242 381
rect 90 341 242 347
rect 422 381 574 387
rect 422 347 434 381
rect 562 347 574 381
rect 422 341 574 347
rect -630 297 -584 309
rect -630 121 -624 297
rect -590 121 -584 297
rect -630 109 -584 121
rect -412 297 -366 309
rect -412 121 -406 297
rect -372 121 -366 297
rect -412 109 -366 121
rect -298 297 -252 309
rect -298 121 -292 297
rect -258 121 -252 297
rect -298 109 -252 121
rect -80 297 -34 309
rect -80 121 -74 297
rect -40 121 -34 297
rect -80 109 -34 121
rect 34 297 80 309
rect 34 121 40 297
rect 74 121 80 297
rect 34 109 80 121
rect 252 297 298 309
rect 252 121 258 297
rect 292 121 298 297
rect 252 109 298 121
rect 366 297 412 309
rect 366 121 372 297
rect 406 121 412 297
rect 366 109 412 121
rect 584 297 630 309
rect 584 121 590 297
rect 624 121 630 297
rect 584 109 630 121
rect -574 71 -422 77
rect -574 37 -562 71
rect -434 37 -422 71
rect -574 31 -422 37
rect -242 71 -90 77
rect -242 37 -230 71
rect -102 37 -90 71
rect -242 31 -90 37
rect 90 71 242 77
rect 90 37 102 71
rect 230 37 242 71
rect 90 31 242 37
rect 422 71 574 77
rect 422 37 434 71
rect 562 37 574 71
rect 422 31 574 37
rect -574 -37 -422 -31
rect -574 -71 -562 -37
rect -434 -71 -422 -37
rect -574 -77 -422 -71
rect -242 -37 -90 -31
rect -242 -71 -230 -37
rect -102 -71 -90 -37
rect -242 -77 -90 -71
rect 90 -37 242 -31
rect 90 -71 102 -37
rect 230 -71 242 -37
rect 90 -77 242 -71
rect 422 -37 574 -31
rect 422 -71 434 -37
rect 562 -71 574 -37
rect 422 -77 574 -71
rect -630 -121 -584 -109
rect -630 -297 -624 -121
rect -590 -297 -584 -121
rect -630 -309 -584 -297
rect -412 -121 -366 -109
rect -412 -297 -406 -121
rect -372 -297 -366 -121
rect -412 -309 -366 -297
rect -298 -121 -252 -109
rect -298 -297 -292 -121
rect -258 -297 -252 -121
rect -298 -309 -252 -297
rect -80 -121 -34 -109
rect -80 -297 -74 -121
rect -40 -297 -34 -121
rect -80 -309 -34 -297
rect 34 -121 80 -109
rect 34 -297 40 -121
rect 74 -297 80 -121
rect 34 -309 80 -297
rect 252 -121 298 -109
rect 252 -297 258 -121
rect 292 -297 298 -121
rect 252 -309 298 -297
rect 366 -121 412 -109
rect 366 -297 372 -121
rect 406 -297 412 -121
rect 366 -309 412 -297
rect 584 -121 630 -109
rect 584 -297 590 -121
rect 624 -297 630 -121
rect 584 -309 630 -297
rect -574 -347 -422 -341
rect -574 -381 -562 -347
rect -434 -381 -422 -347
rect -574 -387 -422 -381
rect -242 -347 -90 -341
rect -242 -381 -230 -347
rect -102 -381 -90 -347
rect -242 -387 -90 -381
rect 90 -347 242 -341
rect 90 -381 102 -347
rect 230 -381 242 -347
rect 90 -387 242 -381
rect 422 -347 574 -341
rect 422 -381 434 -347
rect 562 -381 574 -347
rect 422 -387 574 -381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
