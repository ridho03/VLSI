magic
tech sky130A
magscale 1 2
timestamp 1729184360
<< pwell >>
rect -425 -348 425 348
<< nmos >>
rect -229 -200 -29 200
rect 29 -200 229 200
<< ndiff >>
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
<< ndiffc >>
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
<< psubdiff >>
rect -389 278 -293 312
rect 293 278 389 312
rect -389 216 -355 278
rect 355 216 389 278
rect -389 -278 -355 -216
rect 355 -278 389 -216
rect -389 -312 -293 -278
rect 293 -312 389 -278
<< psubdiffcont >>
rect -293 278 293 312
rect -389 -216 -355 216
rect 355 -216 389 216
rect -293 -312 293 -278
<< poly >>
rect -229 200 -29 226
rect 29 200 229 226
rect -229 -226 -29 -200
rect 29 -226 229 -200
<< locali >>
rect -389 278 -293 312
rect 293 278 389 312
rect -389 216 -355 278
rect 355 216 389 278
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect -389 -278 -355 -216
rect 355 -278 389 -216
rect -389 -312 -293 -278
rect 293 -312 389 -278
<< viali >>
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
<< metal1 >>
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
<< properties >>
string FIXED_BBOX -372 -295 372 295
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
