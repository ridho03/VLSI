magic
tech sky130A
magscale 1 2
timestamp 1729317316
<< psubdiff >>
rect -1070 4424 -1010 4458
rect 2445 4424 2505 4458
rect -1070 4398 -1036 4424
rect -1070 1079 -1036 1105
rect 2471 4398 2505 4424
rect 2471 1079 2505 1105
rect -1070 1045 -1010 1079
rect 2445 1045 2505 1079
<< psubdiffcont >>
rect -1010 4424 2445 4458
rect -1070 1105 -1036 4398
rect 2471 1105 2505 4398
rect -1010 1045 2445 1079
<< locali >>
rect -1070 4424 -1010 4458
rect 2445 4424 2505 4458
rect -1070 4398 -1036 4424
rect -1070 1079 -1036 1105
rect 2471 4398 2505 4424
rect 2471 1079 2505 1105
rect -1070 1045 -1010 1079
rect 2445 1045 2505 1079
<< metal1 >>
rect 726 4368 1610 4408
rect 726 3870 766 4368
rect 1570 4247 1610 4368
rect 978 4030 988 4082
rect 1040 4030 1050 4082
rect -149 3869 766 3870
rect -182 3835 766 3869
rect -149 3830 766 3835
rect 2130 3317 2194 3324
rect 985 3265 995 3317
rect 1047 3265 1057 3317
rect 2130 3265 2137 3317
rect 2189 3265 2194 3317
rect 2130 3259 2194 3265
rect 2355 3315 2407 3321
rect 2355 3257 2407 3263
rect -182 3134 74 3168
rect 40 2840 74 3134
rect 492 3121 498 3173
rect 550 3164 556 3173
rect 550 3130 957 3164
rect 550 3121 556 3130
rect 2361 3062 2401 3257
rect 2248 3022 2401 3062
rect 1279 2911 1285 2963
rect 1337 2911 1343 2963
rect 40 2806 1074 2840
rect -4 2739 232 2774
rect -4 1942 31 2739
rect 197 2478 232 2739
rect 1040 2474 1074 2806
rect 1294 2033 1328 2911
rect 2248 2876 2297 3022
rect 1294 1999 1422 2033
rect -181 1908 31 1942
<< via1 >>
rect 988 4030 1040 4082
rect 995 3265 1047 3317
rect 2137 3265 2189 3317
rect 2355 3263 2407 3315
rect 498 3121 550 3173
rect 1285 2911 1337 2963
<< metal2 >>
rect 988 4082 1040 4092
rect 988 4020 1040 4030
rect 732 3591 741 3651
rect 801 3638 810 3651
rect 801 3604 949 3638
rect 801 3591 810 3604
rect 481 3261 490 3321
rect 550 3317 559 3321
rect 995 3317 1047 3327
rect 550 3265 995 3317
rect 550 3261 559 3265
rect 995 3255 1047 3265
rect 2130 3317 2194 3324
rect 2130 3265 2137 3317
rect 2189 3315 2365 3317
rect 2189 3265 2355 3315
rect 2130 3259 2194 3265
rect 2349 3263 2355 3265
rect 2407 3263 2413 3315
rect 498 3173 550 3179
rect 498 3115 550 3121
rect 1088 2907 1097 2967
rect 1157 2954 1166 2967
rect 1285 2963 1337 2969
rect 1157 2920 1285 2954
rect 1157 2907 1166 2920
rect 1285 2905 1337 2911
rect 1258 2816 1328 2825
rect 1258 2708 1328 2746
rect 1258 2656 1558 2708
<< via2 >>
rect 741 3591 801 3651
rect 490 3261 550 3321
rect 1097 2907 1157 2967
rect 1258 2746 1328 2816
<< metal3 >>
rect 706 3651 822 3684
rect 706 3591 741 3651
rect 801 3591 822 3651
rect 706 3568 822 3591
rect 485 3321 555 3326
rect 299 3261 490 3321
rect 550 3261 555 3321
rect 299 3251 369 3261
rect 485 3256 555 3261
rect -194 3191 369 3251
rect 299 3072 369 3191
rect 299 3004 300 3072
rect 368 3004 369 3072
rect 299 3003 369 3004
rect 1215 3003 1221 3073
rect 1291 3003 1328 3073
rect 300 2998 368 3003
rect 1092 2967 1162 2972
rect 513 2907 1097 2967
rect 1157 2907 1162 2967
rect 513 2728 597 2907
rect 1092 2902 1162 2907
rect 684 2838 745 2840
rect 683 2832 747 2838
rect 1258 2821 1328 3003
rect 683 2762 747 2768
rect 1253 2816 1333 2821
rect 684 2404 745 2762
rect 1253 2746 1258 2816
rect 1328 2746 1333 2816
rect 1253 2741 1333 2746
<< via3 >>
rect 300 3004 368 3072
rect 1221 3003 1291 3073
rect 683 2768 747 2832
<< metal4 >>
rect 1220 3073 1292 3074
rect 299 3072 1221 3073
rect 299 3004 300 3072
rect 368 3004 1221 3072
rect 299 3003 1221 3004
rect 1291 3003 1292 3073
rect 1220 3002 1292 3003
rect 652 2832 772 2858
rect 652 2768 683 2832
rect 747 2768 772 2832
rect 652 2745 772 2768
use lnmos  lnmos_0
timestamp 1729242596
transform 0 -1 2305 1 0 1439
box -306 -130 1578 929
use lpmos  lpmos_0
timestamp 1729250664
transform 1 0 -693 0 1 3229
box 1513 -185 3054 1089
use nmoscs  nmoscs_0
timestamp 1729218614
transform 1 0 -2739 0 1 1178
box 2801 -71 3980 1550
use pmoscs  pmoscs_0
timestamp 1729158256
transform 1 0 -778 0 1 1055
box -232 53 767 2922
<< labels >>
flabel metal1 299 3855 299 3855 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal3 547 2929 547 2929 0 FreeSans 1600 0 0 0 GND
port 1 nsew
flabel metal3 330 3202 330 3202 0 FreeSans 1600 0 0 0 OUT
port 2 nsew
flabel via3 722 2786 722 2786 0 FreeSans 1600 0 0 0 RS
port 3 nsew
flabel metal1 617 3147 617 3147 0 FreeSans 1600 0 0 0 VIN
port 4 nsew
flabel via2 757 3627 757 3627 0 FreeSans 1600 0 0 0 VIP
port 5 nsew
<< end >>
