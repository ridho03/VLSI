magic
tech sky130A
magscale 1 2
timestamp 1729241487
<< nmos >>
rect -80 -131 80 69
<< ndiff >>
rect -138 57 -80 69
rect -138 -119 -126 57
rect -92 -119 -80 57
rect -138 -131 -80 -119
rect 80 57 138 69
rect 80 -119 92 57
rect 126 -119 138 57
rect 80 -131 138 -119
<< ndiffc >>
rect -126 -119 -92 57
rect 92 -119 126 57
<< poly >>
rect -80 141 80 157
rect -80 107 -64 141
rect 64 107 80 141
rect -80 69 80 107
rect -80 -157 80 -131
<< polycont >>
rect -64 107 64 141
<< locali >>
rect -80 107 -64 141
rect 64 107 80 141
rect -126 57 -92 73
rect -126 -135 -92 -119
rect 92 57 126 73
rect 92 -135 126 -119
<< viali >>
rect -45 107 45 141
rect -126 -119 -92 57
rect 92 -119 126 57
<< metal1 >>
rect -57 141 57 147
rect -57 107 -45 141
rect 45 107 57 141
rect -57 101 57 107
rect -132 57 -86 69
rect -132 -119 -126 57
rect -92 -119 -86 57
rect -132 -131 -86 -119
rect 86 57 132 69
rect 86 -119 92 57
rect 126 -119 132 57
rect 86 -131 132 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
