magic
tech sky130A
magscale 1 2
timestamp 1729242596
<< pwell >>
rect -306 -112 1578 916
<< psubdiff >>
rect -306 882 -246 916
rect 1518 882 1578 916
rect -306 856 -272 882
rect 1544 856 1578 882
rect -306 -78 -272 -52
rect 1544 -78 1578 -52
rect -306 -112 -246 -78
rect 1518 -112 1578 -78
<< psubdiffcont >>
rect -246 882 1518 916
rect -306 -52 -272 856
rect 1544 -52 1578 856
rect -246 -112 1518 -78
<< poly >>
rect -160 778 0 794
rect -160 744 -144 778
rect -16 744 0 778
rect -160 718 0 744
rect 1272 778 1432 794
rect 1272 744 1288 778
rect 1416 744 1432 778
rect 1272 717 1432 744
rect 58 376 1214 418
rect -160 50 0 77
rect -160 16 -144 50
rect -16 16 0 50
rect -160 0 0 16
rect 1272 50 1432 77
rect 1272 16 1288 50
rect 1416 16 1432 50
rect 1272 0 1432 16
<< polycont >>
rect -144 744 -16 778
rect 1288 744 1416 778
rect -144 16 -16 50
rect 1288 16 1416 50
<< locali >>
rect -306 882 -246 916
rect 1518 882 1578 916
rect -306 856 -272 882
rect 1544 856 1578 882
rect -160 744 -144 778
rect -16 744 0 778
rect 1272 744 1288 778
rect 1416 744 1432 778
rect -160 16 -144 50
rect -16 16 0 50
rect 1272 16 1288 50
rect 1416 16 1432 50
rect -306 -78 -272 -52
rect 1544 -78 1578 -52
rect -306 -112 -246 -78
rect 1518 -112 1578 -78
<< viali >>
rect 560 916 594 917
rect 560 883 594 916
rect -125 744 -35 778
rect 1307 744 1397 778
rect -125 16 -35 50
rect 1307 16 1397 50
rect 674 -78 710 -77
rect 674 -112 710 -78
rect 674 -113 710 -112
<< metal1 >>
rect 554 917 600 929
rect 554 883 560 917
rect 594 883 600 917
rect 554 874 600 883
rect 224 828 602 874
rect -212 778 0 786
rect -212 744 -125 778
rect -35 744 0 778
rect -212 737 0 744
rect -212 707 -166 737
rect -212 694 56 707
rect 224 697 270 828
rect 556 706 602 828
rect 670 828 1048 874
rect 670 706 716 828
rect 556 694 716 706
rect 1002 698 1048 828
rect 1272 778 1483 786
rect 1272 744 1307 778
rect 1397 744 1483 778
rect 1272 737 1483 744
rect 1438 708 1483 737
rect 1217 694 1485 708
rect -212 518 3 694
rect 55 518 65 694
rect 325 518 335 694
rect 387 518 397 694
rect -212 505 56 518
rect 6 474 52 505
rect 6 428 86 474
rect -212 276 56 289
rect -212 100 3 276
rect 55 100 65 276
rect 325 100 335 276
rect 387 100 397 276
rect -212 87 56 100
rect -212 57 -166 87
rect -212 50 0 57
rect -212 16 -125 50
rect -35 16 0 50
rect -212 8 0 16
rect 224 -24 270 94
rect 557 87 716 694
rect 875 518 885 694
rect 937 518 947 694
rect 1207 518 1217 694
rect 1269 518 1485 694
rect 1217 506 1485 518
rect 1186 320 1266 366
rect 1220 289 1266 320
rect 1216 276 1484 289
rect 875 100 885 276
rect 937 100 947 276
rect 1207 100 1217 276
rect 1269 100 1484 276
rect 557 -24 603 87
rect 224 -70 603 -24
rect 668 -24 716 87
rect 1002 -24 1048 95
rect 1216 87 1484 100
rect 1438 57 1483 87
rect 1272 50 1483 57
rect 1272 16 1307 50
rect 1397 16 1483 50
rect 1272 8 1483 16
rect 668 -70 1048 -24
rect 668 -77 716 -70
rect 668 -113 674 -77
rect 710 -113 716 -77
rect 668 -130 716 -113
<< via1 >>
rect 3 518 55 694
rect 335 518 387 694
rect 3 100 55 276
rect 335 100 387 276
rect 885 518 937 694
rect 1217 518 1269 694
rect 885 100 937 276
rect 1217 100 1269 276
<< metal2 >>
rect 3 794 387 846
rect 3 694 55 794
rect 3 508 55 518
rect 335 694 387 794
rect 885 794 1269 846
rect 885 694 937 794
rect 335 477 387 518
rect 881 518 885 526
rect 1217 694 1269 794
rect 937 518 941 526
rect 335 425 666 477
rect 322 311 331 371
rect 391 311 400 371
rect 614 369 666 425
rect 881 475 941 518
rect 1217 506 1269 518
rect 1226 503 1260 506
rect 881 419 883 475
rect 939 419 941 475
rect 881 417 941 419
rect 883 410 939 417
rect 614 317 937 369
rect 3 276 55 286
rect 3 0 55 100
rect 335 276 387 311
rect 335 0 387 100
rect 3 -52 387 0
rect 885 276 937 317
rect 1226 288 1260 292
rect 885 0 937 100
rect 1217 286 1268 288
rect 1217 276 1269 286
rect 1217 0 1269 100
rect 885 -52 1269 0
<< via2 >>
rect 331 311 391 371
rect 883 419 939 475
<< metal3 >>
rect 878 477 944 480
rect 612 475 944 477
rect 612 419 883 475
rect 939 419 944 475
rect 612 417 944 419
rect 326 371 396 376
rect 612 371 672 417
rect 878 414 944 417
rect 326 311 331 371
rect 391 311 672 371
rect 326 306 396 311
use sky130_fd_pr__nfet_01v8_9C8FNP  sky130_fd_pr__nfet_01v8_9C8FNP_0
timestamp 1729236880
transform 1 0 636 0 1 397
box -636 -397 636 397
use sky130_fd_pr__nfet_01v8_ENL4VF  sky130_fd_pr__nfet_01v8_ENL4VF_0
timestamp 1729241487
transform 1 0 -80 0 1 606
box -138 -126 138 126
use sky130_fd_pr__nfet_01v8_ENL4VF  sky130_fd_pr__nfet_01v8_ENL4VF_1
timestamp 1729241487
transform 1 0 -80 0 1 188
box -138 -126 138 126
use sky130_fd_pr__nfet_01v8_ENL4VF  sky130_fd_pr__nfet_01v8_ENL4VF_3
timestamp 1729241487
transform 1 0 1352 0 1 606
box -138 -126 138 126
use sky130_fd_pr__nfet_01v8_ENL4VF  sky130_fd_pr__nfet_01v8_ENL4VF_4
timestamp 1729241487
transform 1 0 1352 0 1 188
box -138 -126 138 126
<< labels >>
flabel metal1 573 832 573 832 0 FreeSans 1600 0 0 0 gnd
port 0 nsew
flabel metal2 1231 805 1231 805 0 FreeSans 1600 0 0 0 out
port 1 nsew
flabel metal2 29 756 29 756 0 FreeSans 1600 0 0 0 d8
port 2 nsew
<< end >>
