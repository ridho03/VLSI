magic
tech sky130A
magscale 1 2
timestamp 1729250664
<< nwell >>
rect 1513 -185 3054 1089
<< nsubdiff >>
rect 1549 1019 1609 1053
rect 2958 1019 3018 1053
rect 1549 977 1583 1019
rect 2984 977 3018 1019
rect 1549 -115 1583 -89
rect 2984 -115 3018 -89
rect 1549 -149 1609 -115
rect 2958 -149 3018 -115
<< nsubdiffcont >>
rect 1609 1019 2958 1053
rect 1549 -89 1583 977
rect 2984 -89 3018 977
rect 1609 -149 2958 -115
<< poly >>
rect 1674 844 1766 860
rect 1674 810 1690 844
rect 1724 810 1766 844
rect 1674 794 1766 810
rect 1736 785 1766 794
rect 2798 843 2890 859
rect 2798 809 2840 843
rect 2874 809 2890 843
rect 2798 793 2890 809
rect 2798 784 2828 793
rect 1924 465 2096 524
rect 2468 465 2640 522
rect 1924 365 2096 423
rect 2468 365 2640 423
rect 1736 95 1766 104
rect 1674 79 1766 95
rect 1674 45 1690 79
rect 1724 45 1766 79
rect 1674 29 1766 45
rect 2798 95 2828 104
rect 2798 79 2890 95
rect 2798 45 2840 79
rect 2874 45 2890 79
rect 2798 29 2890 45
<< polycont >>
rect 1690 810 1724 844
rect 2840 809 2874 843
rect 1690 45 1724 79
rect 2840 45 2874 79
<< locali >>
rect 1549 1019 1609 1053
rect 2958 1019 3018 1053
rect 1549 977 1583 1019
rect 2984 977 3018 1019
rect 1674 810 1690 844
rect 1724 810 1740 844
rect 1690 746 1724 810
rect 2824 809 2840 843
rect 2874 809 2890 843
rect 2840 734 2874 809
rect 1690 79 1724 141
rect 2840 79 2874 145
rect 1674 45 1690 79
rect 1724 45 1740 79
rect 2824 45 2840 79
rect 2874 45 2890 79
rect 1549 -115 1583 -89
rect 2984 -115 3018 -89
rect 1549 -149 1609 -115
rect 2958 -149 3018 -115
<< viali >>
rect 2264 1019 2302 1053
rect 1690 810 1724 844
rect 2840 809 2874 843
rect 1690 45 1724 79
rect 2840 45 2874 79
<< metal1 >>
rect 2247 1053 2318 1063
rect 2247 1019 2264 1053
rect 2302 1019 2318 1053
rect 2247 1009 2318 1019
rect 1606 947 2964 981
rect 1606 627 1640 947
rect 1936 883 2242 917
rect 1678 844 1736 850
rect 1678 810 1690 844
rect 1724 810 1736 844
rect 1678 804 1736 810
rect 1684 762 1730 804
rect 1836 799 1907 852
rect 1684 750 1821 762
rect 1936 759 1970 883
rect 2109 799 2180 852
rect 2208 762 2242 883
rect 2322 883 2628 917
rect 2322 762 2356 883
rect 2384 801 2455 854
rect 1597 621 1649 627
rect 1597 563 1649 569
rect 1684 574 1769 750
rect 1821 574 1831 750
rect 2031 574 2041 750
rect 2093 574 2103 750
rect 1684 561 1821 574
rect 1840 515 1907 525
rect 1616 481 1907 515
rect 1616 -65 1650 481
rect 1840 472 1907 481
rect 2111 471 2178 524
rect 1683 418 1735 424
rect 1841 409 1908 417
rect 1735 375 1908 409
rect 1683 360 1735 366
rect 1841 364 1908 375
rect 2110 364 2177 417
rect 1684 314 1821 327
rect 1684 138 1769 314
rect 1821 138 1831 314
rect 2031 138 2041 314
rect 2093 138 2103 314
rect 1684 126 1821 138
rect 1684 85 1730 126
rect 1678 79 1736 85
rect 1678 45 1690 79
rect 1724 45 1736 79
rect 1678 39 1736 45
rect 1840 34 1907 87
rect 1936 1 1970 130
rect 2208 126 2356 762
rect 2594 752 2628 883
rect 2660 799 2731 852
rect 2828 843 2886 849
rect 2828 809 2840 843
rect 2874 809 2886 843
rect 2828 803 2886 809
rect 2834 762 2880 803
rect 2743 750 2880 762
rect 2461 574 2471 750
rect 2523 574 2533 750
rect 2733 574 2743 750
rect 2795 574 2880 750
rect 2743 565 2880 574
rect 2389 472 2456 525
rect 2656 515 2723 524
rect 2930 515 2964 947
rect 2656 481 2964 515
rect 2656 471 2723 481
rect 2388 365 2455 418
rect 2658 407 2725 417
rect 2658 373 2963 407
rect 2658 364 2725 373
rect 2743 314 2880 326
rect 2461 138 2471 314
rect 2523 138 2533 314
rect 2733 138 2743 314
rect 2795 138 2880 314
rect 2113 37 2180 90
rect 2208 1 2242 126
rect 1936 -33 2242 1
rect 2322 1 2356 126
rect 2388 38 2455 91
rect 2594 1 2628 132
rect 2743 125 2880 138
rect 2657 35 2724 88
rect 2834 85 2880 125
rect 2828 79 2886 85
rect 2828 45 2840 79
rect 2874 45 2886 79
rect 2828 39 2886 45
rect 2322 -33 2628 1
rect 2929 -65 2963 373
rect 1616 -99 2963 -65
<< via1 >>
rect 1597 569 1649 621
rect 1769 574 1821 750
rect 2041 574 2093 750
rect 1683 366 1735 418
rect 1769 138 1821 314
rect 2041 138 2093 314
rect 2471 574 2523 750
rect 2743 574 2795 750
rect 2471 138 2523 314
rect 2743 138 2795 314
<< metal2 >>
rect 1769 800 2093 852
rect 1769 750 1821 800
rect 1591 569 1597 621
rect 1649 569 1655 621
rect 1606 409 1640 569
rect 1769 564 1821 574
rect 2041 750 2093 800
rect 2041 524 2093 574
rect 2471 800 2795 852
rect 2471 750 2523 800
rect 2471 572 2523 574
rect 2743 750 2795 800
rect 2469 527 2529 572
rect 2743 564 2795 574
rect 2041 472 2305 524
rect 1677 409 1683 418
rect 1606 375 1683 409
rect 1677 366 1683 375
rect 1735 366 1741 418
rect 2028 361 2037 421
rect 2097 361 2106 421
rect 2253 418 2305 472
rect 2469 471 2471 527
rect 2527 471 2529 527
rect 2469 469 2529 471
rect 2471 462 2527 469
rect 2253 366 2523 418
rect 1769 314 1821 324
rect 1769 87 1821 138
rect 2041 314 2093 361
rect 2041 87 2093 138
rect 1769 35 2093 87
rect 2471 314 2523 366
rect 2471 87 2523 138
rect 2743 314 2795 324
rect 2743 87 2795 138
rect 2471 35 2795 87
<< via2 >>
rect 2037 361 2097 421
rect 2471 471 2527 527
<< metal3 >>
rect 2466 529 2532 532
rect 2249 527 2532 529
rect 2249 471 2471 527
rect 2527 471 2532 527
rect 2249 469 2532 471
rect 2032 421 2102 426
rect 2249 421 2309 469
rect 2466 466 2532 469
rect 2032 361 2037 421
rect 2097 361 2309 421
rect 2032 356 2102 361
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729232345
transform 1 0 1751 0 1 226
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729232345
transform 1 0 1751 0 1 662
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729232345
transform 1 0 2813 0 1 662
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729232345
transform 1 0 2813 0 1 226
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_V8A8AU  sky130_fd_pr__pfet_01v8_V8A8AU_0
timestamp 1729243811
transform 1 0 2282 0 1 444
box -552 -418 552 418
<< labels >>
flabel metal2 1795 770 1795 770 0 FreeSans 1280 0 0 0 d6
port 0 nsew
flabel metal1 1824 495 1824 495 0 FreeSans 1280 0 0 0 vin
port 1 nsew
flabel metal1 2771 493 2771 493 0 FreeSans 1280 0 0 0 vip
port 2 nsew
flabel metal2 2769 788 2769 788 0 FreeSans 1280 0 0 0 out
port 3 nsew
flabel metal1 2281 1015 2281 1015 0 FreeSans 1280 0 0 0 vdd
port 4 nsew
<< end >>
